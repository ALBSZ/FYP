clockX = 0
clockY = 0
C = 1
X = 000000000000
Y = 100111000100
P = 000000000000
X_n = 0 0 0 0
Y_n = -276 -20 -4 -4
P_n = 0 0 0 0
X_tmp = 000000000000
Y_tmp = 100111000100
X_increment = 000001000000
Y_increment = 000000000001
X_v = 0
Y_v = -276
P_actual = 0
P_correct = 0
P_C_output = 0
R = 4
D = 3
B = 4
clock_period = 20 ns
